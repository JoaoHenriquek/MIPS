entity PC is
    port (
        in_pc   : in std_logic_vector(15 downto 0);
        out_pc  : in std_logic_vector(15 downto 0);
    );
end PC;

architecture rtl of PC is
begin
    process(out_pc)
    begin
        


begin

end architecture;